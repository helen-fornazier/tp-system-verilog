library verilog;
use verilog.vl_types.all;
entity div_ieee_sv_unit is
end div_ieee_sv_unit;
