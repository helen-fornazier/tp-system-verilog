package float_pack; 
// Ajouter ici les définition des fonctions
// utilisée par votre coprocesseur
endpackage : float_pack
   
