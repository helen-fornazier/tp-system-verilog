import float_pack::*;

module add_ieee(input float op1,
                input float op2,
                output float result
                );
                 
assign result = float_add_sub(1, op1, op2);

endmodule
