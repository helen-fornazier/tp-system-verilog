library verilog;
use verilog.vl_types.all;
entity mult_ieee_sv_unit is
end mult_ieee_sv_unit;
