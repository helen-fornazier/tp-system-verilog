library verilog;
use verilog.vl_types.all;
entity sub_ieee_sv_unit is
end sub_ieee_sv_unit;
