library verilog;
use verilog.vl_types.all;
entity add_ieee_sv_unit is
end add_ieee_sv_unit;
